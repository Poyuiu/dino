module cactus (
        input vsync,
        input clk,
        input rst,
        input [9:0] h_cnt,
        input [9:0] v_cnt,
        input [1:0] state,
        output reg black_cactus
    );
    reg next_black_cactus;

    wire [7:0] rand_num;
    random rand1 (clk, rst, rand_num);

    reg [59:0] ptn0 [57:0];
    reg [59:0] ptn1 [57:0];
    reg [59:0] ptn2 [57:0];
    reg [9:0] cactus_position;
    reg [9:0] next_cactus_position;
    reg [1:0] cactus_type;
    reg [1:0] next_cactus_type;
    reg [9:0] wait_cnt;
    reg [9:0] next_wait_cnt;
    reg [9:0] wait_time;
    reg [9:0] next_wait_time;
    reg last_vsync;
    always @(posedge clk) begin
        if (rst) begin
            cactus_position <= 10'b0;
            last_vsync <= 1'b0;
        end
        else begin
            last_vsync <= vsync;
            if(vsync && !last_vsync && (state != 2'b0 && state != 2'b11)) begin
                if(cactus_position == 10'b0) begin
                    if (wait_cnt == 10'b0) begin
                        wait_time <= (rand_num[3:0]) * 10'd5;//wait time randoms from 0s to 5s (60 frames every second)
                        cactus_type <= (rand_num[4:0]) % 3;//random a cactus type
                        wait_cnt <= 10'b1;
                    end
                    else begin
                        wait_cnt <= wait_cnt + 10'b1;
                        if (wait_cnt >= wait_time) begin//if reached the wait time
                            cactus_position <= 6;//begin to show the cactus
                            wait_cnt <= 10'b0;//make the counter return to zero
                        end
                        else begin
                            cactus_position <= cactus_position;
                        end
                    end
                end
                else begin
                    cactus_position <=
                                    (cactus_position+ 6 )%(10'd640+10'd60);
                end
            end
            else begin
                cactus_position <= cactus_position;
                cactus_type <= cactus_type;
                wait_cnt <= wait_cnt;
                wait_time <= wait_time;
            end
        end
    end

    always @(posedge clk) begin
        if(rst) begin
            black_cactus <= 1'b0;
        end
        else begin
            black_cactus <= next_black_cactus;
        end
    end
    always @(*) begin
        if (v_cnt >= 10'd344 && v_cnt < 10'd402) begin
            if (h_cnt >= (10'd640 > cactus_position ? 10'd640 - cactus_position : 10'd0) && h_cnt < 10'd700 - cactus_position) begin
                //print pattern base on the value of cactus type
                if (cactus_type==0) begin
                    next_black_cactus <= ptn0[v_cnt - 16'd344][h_cnt + cactus_position - 16'd640];
                end
                else if (cactus_type==1) begin
                    next_black_cactus <= ptn1[v_cnt - 16'd344][h_cnt + cactus_position - 16'd640];
                end
                else begin // cactus_type == 2
                    next_black_cactus <= ptn2[v_cnt - 16'd344][h_cnt + cactus_position - 16'd640];
                end
            end
            else begin
                next_black_cactus <= 1'b0;
            end
        end
        else begin
            next_black_cactus <= 1'b0;
        end
    end

    initial begin
        ptn0[0]<=60'b0000000000_0000000000_0000000111_1110000000_0000000000_0000000000;
        ptn0[1]<=60'b0000000000_0000000000_0000001111_1111000000_0000000000_0000000000;
        ptn0[2]<=60'b0000000000_0000000000_0000011111_1111100000_0000000000_0000000000;
        ptn0[3]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[4]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[5]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[6]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[7]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[8]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[9]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[10]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[11]<=60'b0000000000_0000011000_0000111111_1111110000_0000000000_0000000000;
        ptn0[12]<=60'b0000000000_0000111100_0000111111_1111110000_0000000000_0000000000;
        ptn0[13]<=60'b0000000000_0001111110_0000111111_1111110000_0000000000_0000000000;
        ptn0[14]<=60'b0000000000_0011111111_0000111111_1111110000_0011000000_0000000000;
        ptn0[15]<=60'b0000000000_0011111111_0000111111_1111110000_0111100000_0000000000;
        ptn0[16]<=60'b0000000000_0011111111_0000111111_1111110000_1111110000_0000000000;
        ptn0[17]<=60'b0000000000_0011111111_0000111111_1111110000_1111110000_0000000000;
        ptn0[18]<=60'b0000000000_0011111111_0000111111_1111110000_1111110000_0000000000;
        ptn0[19]<=60'b0000000000_0011111111_1111111111_1111110000_1111110000_0000000000;
        ptn0[20]<=60'b0000000000_0011111111_1111111111_1111110000_1111110000_0000000000;
        ptn0[21]<=60'b0000000000_0011111111_1111111111_1111110000_1111110000_0000000000;
        ptn0[22]<=60'b0000000000_0011111111_1111111111_1111110000_1111110000_0000000000;
        ptn0[23]<=60'b0000000000_0011111111_1111111111_1111111111_1111110000_0000000000;
        ptn0[24]<=60'b0000000000_0000111111_1111111111_1111111111_1111110000_0000000000;
        ptn0[25]<=60'b0000000000_0000001111_1111111111_1111111111_1111110000_0000000000;
        ptn0[26]<=60'b0000000000_0000000011_1111111111_1111111111_1111000000_0000000000;
        ptn0[27]<=60'b0000000000_0000000000_1111111111_1111111111_1100000000_0000000000;
        ptn0[28]<=60'b0000000000_0000000000_0000111111_1111111111_0000000000_0000000000;
        ptn0[29]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[30]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[31]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[32]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[33]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[34]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[35]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[36]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[37]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[38]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[39]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[40]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[41]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[42]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[43]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[44]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[45]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[46]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[47]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[48]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[49]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[50]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[51]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[52]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[53]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[54]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[55]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[56]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn0[57]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;


        ptn1[0]<=60'b0000000000_0000000000_0000000111_1110000000_0000000000_0000000000;
        ptn1[1]<=60'b0000000000_0000000000_0000001111_1111000000_0000000000_0000000000;
        ptn1[2]<=60'b0000000000_0000000000_0000011111_1111100000_0000000000_0000000000;
        ptn1[3]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn1[4]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn1[5]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn1[6]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn1[7]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn1[8]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn1[9]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn1[10]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn1[11]<=60'b0000000000_0000011000_0000111111_1111110000_0000000000_0000000000;
        ptn1[12]<=60'b0000000000_0000111100_0000111111_1111110000_0000000000_0000000000;
        ptn1[13]<=60'b0000000000_0001111110_0000111111_1111110000_0000000000_0000000000;
        ptn1[14]<=60'b0000000000_0011111111_0000111111_1111110000_0011000000_0000000000;
        ptn1[15]<=60'b0000000000_0011111111_0000111111_1111110000_0111100000_0000000000;
        ptn1[16]<=60'b0000000000_0011111111_0000111111_1111110000_1111110000_0000000000;
        ptn1[17]<=60'b0000000000_0011111111_0000111111_1111110000_1111110000_0000000000;
        ptn1[18]<=60'b0000000000_0011111111_0000111111_1111110000_1111110000_0000000000;
        ptn1[19]<=60'b0000000000_0011111111_1111111111_1111110000_1111110000_0000000000;
        ptn1[20]<=60'b0000000000_0011111111_1111111111_1111110000_1111110000_0000000000;
        ptn1[21]<=60'b0000000000_0011111111_1111111111_1111110000_1111110000_0000000000;
        ptn1[22]<=60'b0000000000_0011111111_1111111111_1111110000_1111110000_0000000000;
        ptn1[23]<=60'b0000000000_0011111111_1111111111_1111111111_1111110000_0000000000;
        ptn1[24]<=60'b0000000000_0000111111_1111111111_1111111111_1111110000_0000000000;
        ptn1[25]<=60'b0000000000_0000001111_1111111111_1111111111_1111110000_0000000000;
        ptn1[26]<=60'b0000000000_0000000011_1111111111_1111111111_1111000000_0000000000;
        ptn1[27]<=60'b0000000000_0000000000_1111111111_1111111111_1100000000_0000000000;
        ptn1[28]<=60'b0000000000_0000000000_0000111111_1111111111_0000000000_0000000000;
        ptn1[29]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn1[30]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        ptn1[31]<=60'b0000000000_0000000000_0000111111_1111110000_0000000110_0000000000;
        ptn1[32]<=60'b0000000000_0000000000_0000111111_1111110000_0000001111_0000000000;
        ptn1[33]<=60'b0000000000_0000000000_0000111111_1111110000_0000001111_0000000000;
        ptn1[34]<=60'b0000000000_0000000000_0000111111_1111110000_0000001111_0000000000;
        ptn1[35]<=60'b0000000000_0000000000_0000111111_1111110000_0000001111_0000100000;
        ptn1[36]<=60'b0000000000_0000000000_0000111111_1111110000_0000001111_0001110000;
        ptn1[37]<=60'b0000000000_0000000000_0000111111_1111110000_0000001111_0011111000;
        ptn1[38]<=60'b0000000000_0000000000_0000111111_1111110000_0000001111_0011111000;
        ptn1[39]<=60'b0000000000_0000000000_0000111111_1111110000_0000001111_0011111000;
        ptn1[40]<=60'b0000011000_0000000000_0000111111_1111110000_0110001111_0011111000;
        ptn1[41]<=60'b0000111100_0000000000_0000111111_1111110000_1111001111_0011111000;
        ptn1[42]<=60'b0000111100_0000000000_0000111111_1111110000_1111001111_0111110000;
        ptn1[43]<=60'b0000111100_1000000000_0000111111_1111110000_1111001111_1111100000;
        ptn1[44]<=60'b0100111101_1100000000_0000111111_1111110000_1111001111_1111000000;
        ptn1[45]<=60'b1110111101_1100000000_0000111111_1111110000_1111001111_1110000000;
        ptn1[46]<=60'b1110111111_1000000000_0000111111_1111110000_1111001111_1100000000;
        ptn1[47]<=60'b1110111111_0000000000_0000111111_1111110000_1111001111_1000000000;
        ptn1[48]<=60'b1110111110_0000000000_0000111111_1111110000_1111001111_0000000000;
        ptn1[49]<=60'b1110111100_0000000000_0000111111_1111110000_0111101111_0000000000;
        ptn1[50]<=60'b0111111100_0000000000_0000111111_1111110000_0011111111_0000000000;
        ptn1[51]<=60'b0011111100_0000000000_0000111111_1111110000_0001111111_0000000000;
        ptn1[52]<=60'b0001111100_0000000000_0000111111_1111110000_0000111111_0000000000;
        ptn1[53]<=60'b0000111100_0000000000_0000111111_1111110000_0000011111_0000000000;
        ptn1[54]<=60'b0000111100_0000000000_0000111111_1111110000_0000001111_0000000000;
        ptn1[55]<=60'b0000111100_0000000000_0000111111_1111110000_0000001111_0000000000;
        ptn1[56]<=60'b0000111100_0000000000_0000111111_1111110000_0000001111_0000000000;
        ptn1[57]<=60'b0000111100_0000000000_0000111111_1111110000_0000001111_0000000000;

        ptn2[0]<=60'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        ptn2[1]<=60'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        ptn2[2]<=60'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        ptn2[3]<=60'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        ptn2[4]<=60'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        ptn2[5]<=60'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        ptn2[6]<=60'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        ptn2[7]<=60'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        ptn2[8]<=60'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        ptn2[9]<=60'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        ptn2[10]<=60'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        ptn2[11]<=60'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        ptn2[12]<=60'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        ptn2[13]<=60'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        ptn2[14]<=60'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        ptn2[15]<=60'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        ptn2[16]<=60'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        ptn2[17]<=60'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        ptn2[18]<=60'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        ptn2[19]<=60'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        ptn2[20]<=60'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        ptn2[21]<=60'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        ptn2[22]<=60'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        ptn2[23]<=60'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        ptn2[24]<=60'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        ptn2[25]<=60'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        ptn2[26]<=60'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        ptn2[27]<=60'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        ptn2[28]<=60'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        ptn2[29]<=60'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        ptn2[30]<=60'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        ptn2[31]<=60'b0000000000_0000000000_0000000001_1000000000_0000000000_0000000000;
        ptn2[32]<=60'b0000000000_0000000000_0000000011_1100000000_0000000000_0000000000;
        ptn2[33]<=60'b0000000000_0000000000_0000000111_1110000000_0000000000_0000000000;
        ptn2[34]<=60'b0000000000_0000000000_0000000111_1110000000_0000000000_0000000000;
        ptn2[35]<=60'b0000000000_0000000000_0000000111_1110000000_0000000000_0000000000;
        ptn2[36]<=60'b0000000000_0000000000_0000000111_1110000000_0000000000_0000000000;
        ptn2[37]<=60'b0000000000_0000000000_0000000111_1110000000_0000000000_0000000000;
        ptn2[38]<=60'b0000000000_0000000000_0000000111_1110000000_0000000000_0000000000;
        ptn2[39]<=60'b0000000000_0000000000_0000000111_1110000000_0000000000_0000000000;
        ptn2[40]<=60'b0000000000_0000000000_0001000111_1110000000_0000000000_0000000000;
        ptn2[41]<=60'b0000000000_0000000000_0011100111_1110000000_0000000000_0000000000;
        ptn2[42]<=60'b0000000000_0000000000_0011100111_1110000000_0000000000_0000000000;
        ptn2[43]<=60'b0000000000_0000000000_0011100111_1110000000_0000000000_0000000000;
        ptn2[44]<=60'b0000000000_0000000000_0011100111_1110001000_0000000000_0000000000;
        ptn2[45]<=60'b0000000000_0000000000_0011100111_1110011100_0000000000_0000000000;
        ptn2[46]<=60'b0000000000_0000000000_0011111111_1110011100_0000000000_0000000000;
        ptn2[47]<=60'b0000000000_0000000000_0001111111_1110011100_0000000000_0000000000;
        ptn2[48]<=60'b0000000000_0000000000_0000111111_1111111100_0000000000_0000000000;
        ptn2[49]<=60'b0000000000_0000000000_0000011111_1111111000_0000000000_0000000000;
        ptn2[50]<=60'b0000000000_0000000000_0000001111_1111110000_0000000000_0000000000;
        ptn2[51]<=60'b0000000000_0000000000_0000000111_1111100000_0000000000_0000000000;
        ptn2[52]<=60'b0000000000_0000000000_0000000111_1111000000_0000000000_0000000000;
        ptn2[53]<=60'b0000000000_0000000000_0000000111_1110000000_0000000000_0000000000;
        ptn2[54]<=60'b0000000000_0000000000_0000000111_1110000000_0000000000_0000000000;
        ptn2[55]<=60'b0000000000_0000000000_0000000111_1110000000_0000000000_0000000000;
        ptn2[56]<=60'b0000000000_0000000000_0000000111_1110000000_0000000000_0000000000;
        ptn2[57]<=60'b0000000000_0000000000_0000000111_1110000000_0000000000_0000000000;
    end
endmodule
