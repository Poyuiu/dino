module ground (
        input [9:0] h_cnt,
        input [9:0] v_cnt,
        input vsync,
        input clk,
        input [1:0] state,
        input rst,
        output reg black_ground
    );

    reg last_vsync;
    reg [159:0] pattern [7:0];
    initial begin
        pattern[0]<=160'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111;
        pattern[1]<=160'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        pattern[2]<=160'b0000000000_0111000000_0000000000_0000000011_1000000000_0000000000_0000000000_0000000000_0000000110_0000000000_0000000000_0111000000_0000000000_0000000000_0000000000_0000000000;
        pattern[3]<=160'b0000000000_0000000000_0000000000_0000000000_0000110000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000111000_0000000000_0000000000_0000000000;
        pattern[4]<=160'b0000000000_0100000000_0000000000_0000110000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0011000000;
        pattern[5]<=160'b0000000000_0000000000_0000011100_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0011110000_0000000000_0000000000_0000000000_0000000000_0000000000;
        pattern[6]<=160'b0000000010_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0011000000_0000000000_0000000000_0000000000_0000000000_0000000000_1110000000_0000000000_0000000000;
        pattern[7]<=160'b0000000000_0111000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000001000;
    end
    reg [9:0] ground_position;

    always @(posedge clk) begin
        if (rst) begin
            ground_position <= 10'b0;
            last_vsync <= 1'b0;
        end
        else begin
            last_vsync <= vsync;
            if(vsync && !last_vsync && state != 2'b0)
                ground_position<=(ground_position+6)%10'd160;//move the ground
            else
                ground_position <= ground_position;
        end
    end
    reg next_black_ground;
    always @(posedge clk) begin
        if(rst) begin
            black_ground <= 1'b0;
        end
        else begin
            black_ground <= next_black_ground;
        end
    end
    always @(*) begin
        if(v_cnt < 400)
            next_black_ground = 1'b0;
        else if(v_cnt < 408) begin
            next_black_ground =
                (pattern[v_cnt-10'd400][(h_cnt+ground_position)%10'd160] == 1)
                ? 1'b1 : 1'b0;
        end
        else if(v_cnt < 480)
            next_black_ground = 1'b0;
        else
            next_black_ground = 1'b0;
    end
endmodule
