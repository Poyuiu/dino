module jump (
        input clk, //clock signal
        input jump_op, // jump signal for player
        input Q_jump, // jump signal for q learn
        input rst, // reset signal
        input [9:0] h_cnt, // like x coordinate on screen
        input [9:0] v_cnt, // like y coordinate on screen
        input [1:0] state, // game state
        input new_frame, // game clock
        output reg black_dino, // pixel
        output reg success_jump, // send back to bot(Qlearn), let it check if jump success
        output reg jumping // send back to bot(Qlearn), let it setect the action
    );

    // game states
    parameter INITIAL = 2'b00;
    parameter PLAY = 2'b01;
    parameter Q_LEARNING = 2'b10;
    parameter DEAD = 2'b11;

    // how much time process after jumping
    reg [11:0] jump_time;
    // use jump_time to compute appropriate height the dino should be
    wire [11:0] height;
    // the dino appearance
    reg [0:82] body_run [0:73];
    reg [0:82] body_stop [0:73];
    reg [0:82] feet_stop [0:13];
    reg [0:82] feet_run_a [0:13];
    reg [0:82] feet_run_b [0:13];
    //determine the speed the dino's foot alternate
    reg [3:0] counter;

    //height is only associated with the value of jump_time
    assign height = (jump_time*12'd40 - jump_time*jump_time) / 2'd2;

    //for every frame
    always @(posedge clk) begin
        if(rst) begin
            counter <= 4'b0;
            jumping <= 1'b0;
            jump_time <= 12'b0;
        end
        else begin
            if(new_frame) begin // game clock update every parameter in the game
                counter <= counter+4'b1; // used for running foot
                case (state)
                    INITIAL: begin
                        // initial state
                        success_jump <= 1'b0;
                        if(jump_op) begin // set if jumping
                            jump_time <= 12'b0;
                            jumping <= 1'b1;
                        end
                        else begin
                            jump_time <= 12'b0;
                            jumping <= 1'b0;
                        end
                    end
                    PLAY: begin
                        // playing
                        success_jump <= 1'b0;
                        if (jump_op && jumping==1'b0) begin //begin to jump
                            jumping <= 1'b1;
                            jump_time <= jump_time;
                        end
                        else if (jumping) begin // during jumping
                            if (jump_time >= 12'd40) begin // reset jump operation
                                jump_time <= 12'b0;
                                jumping <= 1'b0;
                            end
                            else begin
                                jumping <= jumping;
                                jump_time <= jump_time+12'b1; // add jump_time
                            end
                        end
                        else begin // nothing -> keep
                            jumping <= jumping;
                            jump_time <= jump_time;
                        end
                    end
                    Q_LEARNING: begin // Q learning
                        if (Q_jump && jumping==1'b0) begin //begin to jump
                            jumping <= 1'b1;
                            // set for bot, the timing dino jump
                            // just one game clock cycle
                            success_jump <= 1'b1;
                            jump_time <= jump_time;
                        end
                        else if (jumping) begin
                            success_jump <= 1'b0; // set to 0
                            if (jump_time >= 12'd40) begin // reset jump operation
                                jump_time <= 12'b0;
                                jumping <= 1'b0;
                            end
                            else begin
                                jumping <= jumping;
                                jump_time <= jump_time+12'b1; // add jump_time
                            end
                        end
                        else begin
                            success_jump <= 1'b0; // set to 0
                            jumping <= jumping;
                            jump_time <= jump_time;
                        end
                    end
                    default: begin
                        // DEAD state
                        success_jump <= 1'b0;
                        jump_time <= jump_time;
                        jumping <= jumping;
                    end
                endcase
            end
            else begin // when game clock isn't triggered -> keep
                counter <= counter;
                success_jump <= 1'b0;
                jumping <= jumping;
                jump_time <= jump_time;
            end
        end
    end
    // check the coordinate to set the pixel signal
    always @(posedge clk) begin
        if(rst) begin
            black_dino <= 1'b0;
        end
        else begin
            // the possible position the dino's body appears
            if (v_cnt >= 10'd402 - height - 10'd88 && v_cnt < 10'd402 - height -10'd14 && h_cnt>=10'd80 && h_cnt<10'd162) begin
                if (state == 2'b11) begin // if it stops
                    black_dino <= body_stop[v_cnt+height-10'd314][h_cnt-10'd80];
                end
                else  begin // if running
                    black_dino <= body_run[v_cnt+height-10'd314][h_cnt-10'd80];
                end

            end
            else begin
                black_dino <= 1'b0;
            end
            // the possible position the dino's feet appears
            if (v_cnt >= 10'd402 - height - 10'd14 && v_cnt < 10'd402 - height && h_cnt>=10'd80 && h_cnt<10'd162) begin
                if ((state != 2'b0 && state != 2'b11) && height==0) begin
                    // moving feet
                    if (counter[3]) begin
                        black_dino <= feet_run_a[v_cnt+height-10'd388][h_cnt-10'd80];
                    end
                    else begin
                        black_dino <= feet_run_b[v_cnt+height-10'd388][h_cnt-10'd80];
                    end
                end
                else begin
                    // stopped feet
                    black_dino <= feet_stop[v_cnt+height-10'd388][h_cnt-10'd80];
                end

            end
        end
    end
    // initial every status dino by always and rst signal
    // reg array reference: https://github.com/awmleer/dinosaur
    always @(posedge clk) begin
        if(rst) begin
            body_run[0]<=82'b0000000000_0000000000_0000000000_0000000000_0000000011_1111111111_1111111111_1111111100_00;
            body_run[1]<=82'b0000000000_0000000000_0000000000_0000000000_0000000011_1111111111_1111111111_1111111100_00;
            body_run[2]<=82'b0000000000_0000000000_0000000000_0000000000_0000000011_1111111111_1111111111_1111111100_00;
            body_run[3]<=82'b0000000000_0000000000_0000000000_0000000000_0000000011_1111111111_1111111111_1111111100_00;
            body_run[4]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
            body_run[5]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
            body_run[6]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
            body_run[7]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
            body_run[8]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1100011111_1111111111_1111111111_11;
            body_run[9]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1100011111_1111111111_1111111111_11;
            body_run[10]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1100011111_1111111111_1111111111_11;
            body_run[11]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
            body_run[12]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
            body_run[13]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
            body_run[14]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
            body_run[15]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
            body_run[16]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
            body_run[17]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
            body_run[18]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
            body_run[19]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
            body_run[20]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
            body_run[21]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
            body_run[22]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
            body_run[23]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1110000000_0000000000_00;
            body_run[24]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1110000000_0000000000_00;
            body_run[25]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1110000000_0000000000_00;
            body_run[26]<=82'b1111000000_0000000000_0000000000_0000000000_1111111111_1111111111_1111111111_1111111100_00;
            body_run[27]<=82'b1111000000_0000000000_0000000000_0000000000_1111111111_1111111111_1111111111_1111111100_00;
            body_run[28]<=82'b1111000000_0000000000_0000000000_0000001111_1111111111_1111110000_0000000000_0000000000_00;
            body_run[29]<=82'b1111000000_0000000000_0000000000_0000001111_1111111111_1111110000_0000000000_0000000000_00;
            body_run[30]<=82'b1111000000_0000000000_0000000000_0000111111_1111111111_1111110000_0000000000_0000000000_00;
            body_run[31]<=82'b1111000000_0000000000_0000000000_0000111111_1111111111_1111110000_0000000000_0000000000_00;
            body_run[32]<=82'b1111110000_0000000000_0000000000_0011111111_1111111111_1111110000_0000000000_0000000000_00;
            body_run[33]<=82'b1111110000_0000000000_0000000000_0011111111_1111111111_1111110000_0000000000_0000000000_00;
            body_run[34]<=82'b1111111100_0000000000_0000000000_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_run[35]<=82'b1111111100_0000000000_0000000000_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_run[36]<=82'b1111111111_0000000000_0000001111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_run[37]<=82'b1111111111_0000000000_0000001111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_run[38]<=82'b1111111111_1100000000_0000111111_1111111111_1111111111_1111111111_1111000000_0000000000_00;
            body_run[39]<=82'b1111111111_1100000000_0000111111_1111111111_1111111111_1111111111_1111000000_0000000000_00;
            body_run[40]<=82'b1111111111_1111000000_1111111111_1111111111_1111111111_1111111111_1111000000_0000000000_00;
            body_run[41]<=82'b1111111111_1111000000_1111111111_1111111111_1111111111_1111111111_1111000000_0000000000_00;
            body_run[42]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_1111000000_0000000000_00;
            body_run[43]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_1111000000_0000000000_00;
            body_run[44]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_1111000000_0000000000_00;
            body_run[45]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_1111000000_0000000000_00;
            body_run[46]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_run[47]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_run[48]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_run[49]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_run[50]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_run[51]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_run[52]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_run[53]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_run[54]<=82'b0011111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_run[55]<=82'b0011111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_run[56]<=82'b0000111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_run[57]<=82'b0000111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_run[58]<=82'b0000001111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_run[59]<=82'b0000001111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_run[60]<=82'b0000000011_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_run[61]<=82'b0000000011_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_run[62]<=82'b0000000000_1111111111_1111111111_1111111111_1111111111_1111000000_0000000000_0000000000_00;
            body_run[63]<=82'b0000000000_1111111111_1111111111_1111111111_1111111111_1111000000_0000000000_0000000000_00;
            body_run[64]<=82'b0000000000_0011111111_1111111111_1111111111_1111111111_1100000000_0000000000_0000000000_00;
            body_run[65]<=82'b0000000000_0011111111_1111111111_1111111111_1111111111_1100000000_0000000000_0000000000_00;
            body_run[66]<=82'b0000000000_0000111111_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000_00;
            body_run[67]<=82'b0000000000_0000111111_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000_00;
            body_run[68]<=82'b0000000000_0000001111_1111111111_1111111111_1111111100_0000000000_0000000000_0000000000_00;
            body_run[69]<=82'b0000000000_0000001111_1111111111_1111111111_1111111100_0000000000_0000000000_0000000000_00;
            body_run[70]<=82'b0000000000_0000000011_1111111111_1111111111_1111110000_0000000000_0000000000_0000000000_00;
            body_run[71]<=82'b0000000000_0000000011_1111111111_1111111111_1111110000_0000000000_0000000000_0000000000_00;
            body_run[72]<=82'b0000000000_0000000000_1111111111_1111111111_1111000000_0000000000_0000000000_0000000000_00;
            body_run[73]<=82'b0000000000_0000000000_1111111111_1111111111_1111000000_0000000000_0000000000_0000000000_00;


            feet_stop[0]<=82'b0000000000_0000000000_1111111111_1100001111_1111000000_0000000000_0000000000_0000000000_00;
            feet_stop[1]<=82'b0000000000_0000000000_1111111111_1100001111_1111000000_0000000000_0000000000_0000000000_00;
            feet_stop[2]<=82'b0000000000_0000000000_1111111100_0000000000_1111000000_0000000000_0000000000_0000000000_00;
            feet_stop[3]<=82'b0000000000_0000000000_1111111100_0000000000_1111000000_0000000000_0000000000_0000000000_00;
            feet_stop[4]<=82'b0000000000_0000000000_1111111100_0000000000_1111000000_0000000000_0000000000_0000000000_00;
            feet_stop[5]<=82'b0000000000_0000000000_1111110000_0000000000_1111000000_0000000000_0000000000_0000000000_00;
            feet_stop[6]<=82'b0000000000_0000000000_1111000000_0000000000_1111000000_0000000000_0000000000_0000000000_00;
            feet_stop[7]<=82'b0000000000_0000000000_1111000000_0000000000_1111000000_0000000000_0000000000_0000000000_00;
            feet_stop[8]<=82'b0000000000_0000000000_1111000000_0000000000_1111000000_0000000000_0000000000_0000000000_00;
            feet_stop[9]<=82'b0000000000_0000000000_1111000000_0000000000_1111000000_0000000000_0000000000_0000000000_00;
            feet_stop[10]<=82'b0000000000_0000000000_1111111100_0000000000_1111111100_0000000000_0000000000_0000000000_00;
            feet_stop[11]<=82'b0000000000_0000000000_1111111100_0000000000_1111111100_0000000000_0000000000_0000000000_00;
            feet_stop[12]<=82'b0000000000_0000000000_1111111100_0000000000_1111111100_0000000000_0000000000_0000000000_00;
            feet_stop[13]<=82'b0000000000_0000000000_1111111100_0000000000_1111111100_0000000000_0000000000_0000000000_00;


            feet_run_a[0]<=82'b0000000000_0000000000_1111111100_0000001111_1111000000_0000000000_0000000000_0000000000_00;
            feet_run_a[1]<=82'b0000000000_0000000000_1111111100_0000001111_1111000000_0000000000_0000000000_0000000000_00;
            feet_run_a[2]<=82'b0000000000_0000000000_1111111100_0000000000_1111000000_0000000000_0000000000_0000000000_00;
            feet_run_a[3]<=82'b0000000000_0000000000_0011111111_1111000000_1111000000_0000000000_0000000000_0000000000_00;
            feet_run_a[4]<=82'b0000000000_0000000000_0011111111_1111000000_1111000000_0000000000_0000000000_0000000000_00;
            feet_run_a[5]<=82'b0000000000_0000000000_0000000000_0000000000_1111000000_0000000000_0000000000_0000000000_00;
            feet_run_a[6]<=82'b0000000000_0000000000_0000000000_0000000000_1111000000_0000000000_0000000000_0000000000_00;
            feet_run_a[7]<=82'b0000000000_0000000000_0000000000_0000000000_1111000000_0000000000_0000000000_0000000000_00;
            feet_run_a[8]<=82'b0000000000_0000000000_0000000000_0000000000_1111000000_0000000000_0000000000_0000000000_00;
            feet_run_a[9]<=82'b0000000000_0000000000_0000000000_0000000000_1111000000_0000000000_0000000000_0000000000_00;
            feet_run_a[10]<=82'b0000000000_0000000000_0000000000_0000000000_1111111100_0000000000_0000000000_0000000000_00;
            feet_run_a[11]<=82'b0000000000_0000000000_0000000000_0000000000_1111111100_0000000000_0000000000_0000000000_00;
            feet_run_a[12]<=82'b0000000000_0000000000_0000000000_0000000000_1111111100_0000000000_0000000000_0000000000_00;
            feet_run_a[13]<=82'b0000000000_0000000000_0000000000_0000000000_1111111100_0000000000_0000000000_0000000000_00;


            feet_run_b[0]<=82'b0000000000_0000000000_1111111111_1100000000_1111000000_0000000000_0000000000_0000000000_00;
            feet_run_b[1]<=82'b0000000000_0000000000_1111111111_1100000000_1111000000_0000000000_0000000000_0000000000_00;
            feet_run_b[2]<=82'b0000000000_0000000000_1111111100_0000000000_1111111111_0000000000_0000000000_0000000000_00;
            feet_run_b[3]<=82'b0000000000_0000000000_1111111100_0000000000_1111111111_0000000000_0000000000_0000000000_00;
            feet_run_b[4]<=82'b0000000000_0000000000_1111111100_0000000000_0000000000_0000000000_0000000000_0000000000_00;
            feet_run_b[5]<=82'b0000000000_0000000000_1111110000_0000000000_0000000000_0000000000_0000000000_0000000000_00;
            feet_run_b[6]<=82'b0000000000_0000000000_1111000000_0000000000_0000000000_0000000000_0000000000_0000000000_00;
            feet_run_b[7]<=82'b0000000000_0000000000_1111000000_0000000000_0000000000_0000000000_0000000000_0000000000_00;
            feet_run_b[8]<=82'b0000000000_0000000000_1111000000_0000000000_0000000000_0000000000_0000000000_0000000000_00;
            feet_run_b[9]<=82'b0000000000_0000000000_1111000000_0000000000_0000000000_0000000000_0000000000_0000000000_00;
            feet_run_b[10]<=82'b0000000000_0000000000_1111111100_0000000000_0000000000_0000000000_0000000000_0000000000_00;
            feet_run_b[11]<=82'b0000000000_0000000000_1111111100_0000000000_0000000000_0000000000_0000000000_0000000000_00;
            feet_run_b[12]<=82'b0000000000_0000000000_1111111100_0000000000_0000000000_0000000000_0000000000_0000000000_00;
            feet_run_b[13]<=82'b0000000000_0000000000_1111111100_0000000000_0000000000_0000000000_0000000000_0000000000_00;



            body_stop[0]<=82'b0000000000_0000000000_0000000000_0000000000_0000000011_1111111111_1111111111_1111111100_00;
            body_stop[1]<=82'b0000000000_0000000000_0000000000_0000000000_0000000011_1111111111_1111111111_1111111100_00;
            body_stop[2]<=82'b0000000000_0000000000_0000000000_0000000000_0000000011_1111111111_1111111111_1111111100_00;
            body_stop[3]<=82'b0000000000_0000000000_0000000000_0000000000_0000000011_1111111111_1111111111_1111111100_00;
            body_stop[4]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
            body_stop[5]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
            body_stop[6]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_0000001111_1111111111_1111111111_11;
            body_stop[7]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_0000001111_1111111111_1111111111_11;
            body_stop[8]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_0011001111_1111111111_1111111111_11;
            body_stop[9]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_0011001111_1111111111_1111111111_11;
            body_stop[10]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_0000001111_1111111111_1111111111_11;
            body_stop[11]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_0000001111_1111111111_1111111111_11;
            body_stop[12]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
            body_stop[13]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
            body_stop[14]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
            body_stop[15]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
            body_stop[16]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
            body_stop[17]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
            body_stop[18]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
            body_stop[19]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
            body_stop[20]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
            body_stop[21]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
            body_stop[22]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
            body_stop[23]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
            body_stop[24]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111100_00;
            body_stop[25]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111100_00;
            body_stop[26]<=82'b1111000000_0000000000_0000000000_0000000000_1111111111_1111111111_1111111111_1111111100_00;
            body_stop[27]<=82'b1111000000_0000000000_0000000000_0000000000_1111111111_1111111111_1111111111_1111111100_00;
            body_stop[28]<=82'b1111000000_0000000000_0000000000_0000001111_1111111111_1111110000_0000000000_0000000000_00;
            body_stop[29]<=82'b1111000000_0000000000_0000000000_0000001111_1111111111_1111110000_0000000000_0000000000_00;
            body_stop[30]<=82'b1111000000_0000000000_0000000000_0000111111_1111111111_1111110000_0000000000_0000000000_00;
            body_stop[31]<=82'b1111000000_0000000000_0000000000_0000111111_1111111111_1111110000_0000000000_0000000000_00;
            body_stop[32]<=82'b1111110000_0000000000_0000000000_0011111111_1111111111_1111110000_0000000000_0000000000_00;
            body_stop[33]<=82'b1111110000_0000000000_0000000000_0011111111_1111111111_1111110000_0000000000_0000000000_00;
            body_stop[34]<=82'b1111111100_0000000000_0000000000_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_stop[35]<=82'b1111111100_0000000000_0000000000_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_stop[36]<=82'b1111111111_0000000000_0000001111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_stop[37]<=82'b1111111111_0000000000_0000001111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_stop[38]<=82'b1111111111_1100000000_0000111111_1111111111_1111111111_1111111111_1111000000_0000000000_00;
            body_stop[39]<=82'b1111111111_1100000000_0000111111_1111111111_1111111111_1111111111_1111000000_0000000000_00;
            body_stop[40]<=82'b1111111111_1111000000_1111111111_1111111111_1111111111_1111111111_1111000000_0000000000_00;
            body_stop[41]<=82'b1111111111_1111000000_1111111111_1111111111_1111111111_1111111111_1111000000_0000000000_00;
            body_stop[42]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_1111000000_0000000000_00;
            body_stop[43]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_1111000000_0000000000_00;
            body_stop[44]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_1111000000_0000000000_00;
            body_stop[45]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_1111000000_0000000000_00;
            body_stop[46]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_stop[47]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_stop[48]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_stop[49]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_stop[50]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_stop[51]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_stop[52]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_stop[53]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_stop[54]<=82'b0011111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_stop[55]<=82'b0011111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_stop[56]<=82'b0000111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_stop[57]<=82'b0000111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_stop[58]<=82'b0000001111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_stop[59]<=82'b0000001111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_stop[60]<=82'b0000000011_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_stop[61]<=82'b0000000011_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
            body_stop[62]<=82'b0000000000_1111111111_1111111111_1111111111_1111111111_1111000000_0000000000_0000000000_00;
            body_stop[63]<=82'b0000000000_1111111111_1111111111_1111111111_1111111111_1111000000_0000000000_0000000000_00;
            body_stop[64]<=82'b0000000000_0011111111_1111111111_1111111111_1111111111_1100000000_0000000000_0000000000_00;
            body_stop[65]<=82'b0000000000_0011111111_1111111111_1111111111_1111111111_1100000000_0000000000_0000000000_00;
            body_stop[66]<=82'b0000000000_0000111111_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000_00;
            body_stop[67]<=82'b0000000000_0000111111_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000_00;
            body_stop[68]<=82'b0000000000_0000001111_1111111111_1111111111_1111111100_0000000000_0000000000_0000000000_00;
            body_stop[69]<=82'b0000000000_0000001111_1111111111_1111111111_1111111100_0000000000_0000000000_0000000000_00;
            body_stop[70]<=82'b0000000000_0000000011_1111111111_1111111111_1111110000_0000000000_0000000000_0000000000_00;
            body_stop[71]<=82'b0000000000_0000000011_1111111111_1111111111_1111110000_0000000000_0000000000_0000000000_00;
            body_stop[72]<=82'b0000000000_0000000000_1111111111_1111111111_1111000000_0000000000_0000000000_0000000000_00;
            body_stop[73]<=82'b0000000000_0000000000_1111111111_1111111111_1111000000_0000000000_0000000000_0000000000_00;
        end
    end
endmodule
